library verilog;
use verilog.vl_types.all;
entity RISC_VDATAPATH_DW01_inc_0 is
    port(
        A               : in     vl_logic_vector(31 downto 0);
        SUM             : out    vl_logic_vector(31 downto 0)
    );
end RISC_VDATAPATH_DW01_inc_0;
